CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 9 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 141 130 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89883e-315 0
0
9 CC 7-Seg~
183 764 135 0 18 19
10 13 12 11 10 9 8 7 18 19
0 0 0 0 0 0 1 2 2
0
0 0 21088 0
6 BLUECC
13 -41 55 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
391 0 0
2
5.89883e-315 5.26354e-315
0
2 +V
167 200 139 0 1 3
0 6
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
5.89883e-315 5.30499e-315
0
6 74LS48
188 662 308 0 14 29
0 5 4 3 2 20 21 7 8 9
10 11 12 13 22
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3421 0 0
2
5.89883e-315 5.32571e-315
0
9 2-In AND~
219 517 94 0 3 22
0 15 4 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8157 0 0
2
5.89883e-315 5.34643e-315
0
9 2-In AND~
219 386 96 0 3 22
0 2 3 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
5.89883e-315 5.3568e-315
0
7 Pulser~
4 82 261 0 10 12
0 23 24 16 25 0 0 5 5 4
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8901 0 0
2
5.89883e-315 5.36716e-315
0
6 74112~
219 580 223 0 7 32
0 6 14 16 14 6 26 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
7361 0 0
2
5.89883e-315 5.37752e-315
0
6 74112~
219 451 224 0 7 32
0 6 15 16 15 6 27 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
4747 0 0
2
5.89883e-315 5.38788e-315
0
6 74112~
219 321 224 0 7 32
0 6 2 16 2 6 28 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
972 0 0
2
5.89883e-315 5.39306e-315
0
6 74112~
219 200 224 0 7 32
0 6 17 16 17 6 29 2
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3472 0 0
2
5.89883e-315 5.39824e-315
0
35
4 0 2 0 0 4224 0 4 0 0 29 3
630 299
237 299
237 188
0 3 3 0 0 12416 0 0 4 26 0 4
349 174
407 174
407 290
630 290
0 2 4 0 0 8320 0 0 4 22 0 4
489 179
546 179
546 281
630 281
7 1 5 0 0 8320 0 8 4 0 0 4
604 187
622 187
622 272
630 272
5 0 6 0 0 12288 0 8 0 0 9 4
580 235
580 239
528 239
528 148
5 0 6 0 0 12288 0 9 0 0 9 4
451 236
451 240
518 240
518 148
5 0 6 0 0 0 0 10 0 0 10 4
321 236
321 240
384 240
384 148
5 0 6 0 0 0 0 11 0 0 11 4
200 236
200 240
259 240
259 148
1 0 6 0 0 8192 0 8 0 0 10 3
580 160
580 148
451 148
1 0 6 0 0 8320 0 9 0 0 11 3
451 161
451 148
321 148
1 1 6 0 0 0 0 10 3 0 0 3
321 161
321 148
200 148
1 1 6 0 0 0 0 3 11 0 0 2
200 148
200 161
7 7 7 0 0 4224 0 2 4 0 0 3
779 171
779 272
694 272
8 6 8 0 0 8320 0 4 2 0 0 3
694 281
773 281
773 171
9 5 9 0 0 8320 0 4 2 0 0 3
694 290
767 290
767 171
10 4 10 0 0 8320 0 4 2 0 0 3
694 299
761 299
761 171
11 3 11 0 0 8320 0 4 2 0 0 3
694 308
755 308
755 171
12 2 12 0 0 8320 0 4 2 0 0 3
694 317
749 317
749 171
13 1 13 0 0 8320 0 4 2 0 0 3
694 326
743 326
743 171
4 0 14 0 0 8192 0 8 0 0 21 3
556 205
542 205
542 186
3 2 14 0 0 8320 0 5 8 0 0 4
538 94
542 94
542 187
556 187
2 7 4 0 0 0 0 5 9 0 0 4
493 103
489 103
489 188
475 188
1 0 15 0 0 4096 0 5 0 0 25 3
493 85
412 85
412 96
0 4 15 0 0 0 0 0 9 25 0 4
412 187
413 187
413 206
427 206
3 2 15 0 0 8320 0 6 9 0 0 4
407 96
412 96
412 188
427 188
2 7 3 0 0 0 0 6 10 0 0 4
362 105
349 105
349 188
345 188
1 0 2 0 0 0 0 6 0 0 28 3
362 87
282 87
282 188
4 0 2 0 0 0 0 10 0 0 29 3
297 206
282 206
282 188
7 2 2 0 0 0 0 11 10 0 0 2
224 188
297 188
3 0 16 0 0 8192 0 8 0 0 31 3
550 196
550 252
418 252
3 0 16 0 0 0 0 9 0 0 32 4
421 197
418 197
418 252
291 252
3 0 16 0 0 8320 0 10 0 0 35 3
291 197
291 252
120 252
1 0 17 0 0 8320 0 1 0 0 34 3
153 130
163 130
163 188
2 4 17 0 0 0 0 11 11 0 0 4
176 188
162 188
162 206
176 206
3 3 16 0 0 0 0 11 7 0 0 4
170 197
120 197
120 252
106 252
1
-32 0 0 0 700 255 0 0 0 3 2 1 18
8 Elephant
0 0 0 12
153 394 491 455
172 402 471 443
12 GALVE, JODIE
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
